module stlb#()();
endmodule