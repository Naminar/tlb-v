module mmu
(
    input translate, // if miss in tlb or significant request
    input [63:0] va,
    input [11:0] pcid
    ouput [63:0] ta
);
    

endmodule